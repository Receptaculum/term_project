`timescale 1ns / 1ps
module decoder(input [3:0] d, output reg [7:0] q);

    always @(*) begin
        case (d)
            4'b0000 : q <= 8'b1111_1100; // 0출력
            4'b0001 : q <= 8'b0110_0000; // 1출력
            4'b0010 : q <= 8'b1101_1010; // 2출력
            4'b0011 : q <= 8'b1111_0010; // 3출력
            4'b0100 : q <= 8'b0110_0110; // 4출력
            4'b0101 : q <= 8'b1011_0110; // 5출력
            4'b0110 : q <= 8'b1011_1110; // 6출력
            4'b0111 : q <= 8'b1110_0100; // 7출력
            4'b1000 : q <= 8'b1111_1110; // 8출력 
            4'b1001 : q <= 8'b1111_0110; // 9출력
        endcase
    end
endmodule